LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY deslocador IS
	PORT(A, B : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		  Dir : IN STD_LOGIC;
		  S : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END deslocador;

ARCHITECTURE arch OF deslocador IS
BEGIN
	PROCESS(A, B, Dir)
	BEGIN
		IF (Dir = '0') THEN
			IF (B = "0000000000000000") THEN
				S <= A;
			ELSIF (B = "0000000000000001") THEN
				S <= A(14 DOWNTO 0) & '0';
			ELSIF (B = "0000000000000010") THEN
				S <= A(13 DOWNTO 0) & "00";
			ELSIF (B = "0000000000000011") THEN
				S <= A(12 DOWNTO 0) & "000";
			ELSIF (B = "0000000000000100") THEN
				S <= A(11 DOWNTO 0) & "0000";
			ELSIF (B = "0000000000000101") THEN
				S <= A(10 DOWNTO 0) & "00000";
			ELSIF (B = "0000000000000110") THEN
				S <= A(9 DOWNTO 0) & "000000";
			ELSIF (B = "0000000000000111") THEN
				S <= A(8 DOWNTO 0) & "0000000";
			ELSIF (B = "0000000000001000") THEN
				S <= A(7 DOWNTO 0) & "00000000";
			ELSIF (B = "0000000000001001") THEN
				S <= A(6 DOWNTO 0) & "000000000";
			ELSIF (B = "0000000000001010") THEN
				S <= A(5 DOWNTO 0) & "0000000000";
			ELSIF (B = "0000000000001011") THEN
				S <= A(4 DOWNTO 0) & "00000000000";
			ELSIF (B = "0000000000001100") THEN
				S <= A(3 DOWNTO 0) & "000000000000";
			ELSIF (B = "0000000000001101") THEN
				S <= A(2 DOWNTO 0) & "0000000000000";
			ELSIF (B = "0000000000001110") THEN
				S <= A(1 DOWNTO 0) & "00000000000000";
			ELSIF (B = "0000000000001111") THEN
				S <= A(0) & "000000000000000";
			ELSE
				S <= "0000000000000000";
			END IF;
		ELSE
			IF (B = "0000000000000000") THEN
				S <= A;
			ELSIF (B = "0000000000000001") THEN
				S <= '0' & A(15 DOWNTO 1);
			ELSIF (B = "0000000000000010") THEN
				S <= "00" & A(15 DOWNTO 2);
			ELSIF (B = "0000000000000011") THEN
				S <= "000" & A(15 DOWNTO 3);
			ELSIF (B = "0000000000000100") THEN
				S <= "0000" & A(15 DOWNTO 4);
			ELSIF (B = "0000000000000101") THEN
				S <= "00000" & A(15 DOWNTO 5);
			ELSIF (B = "0000000000000110") THEN
				S <= "000000" & A(15 DOWNTO 6);
			ELSIF (B = "0000000000000111") THEN
				S <= "0000000" & A(15 DOWNTO 7);
			ELSIF (B = "0000000000001000") THEN
				S <= "00000000" & A(15 DOWNTO 8);
			ELSIF (B = "0000000000001001") THEN
				S <= "000000000" & A(15 DOWNTO 9);
			ELSIF (B = "0000000000001010") THEN
				S <= "0000000000"& A(15 DOWNTO 10);
			ELSIF (B = "0000000000001011") THEN
				S <= "00000000000" & A(15 DOWNTO 11);
			ELSIF (B = "0000000000001100") THEN
				S <= "000000000000" & A(15 DOWNTO 12);
			ELSIF (B = "0000000000001101") THEN
				S <= "0000000000000" & A(15 DOWNTO 13);
			ELSIF (B = "0000000000001110") THEN
				S <= "00000000000000" & A(15 DOWNTO 14);
			ELSIF (B = "0000000000001111") THEN
				S <= "000000000000000" & A(15);
			ELSE
				S <= "0000000000000000";
			END IF;
		END IF;
	END PROCESS;
END;