LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY extensao IS
	PORT(E : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		  S : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END extensao;

ARCHITECTURE arch OF extensao IS
BEGIN
	S <= E(10) & E(10) & E(10) & E(10) & E(10) & E;
END arch;